library verilog;
use verilog.vl_types.all;
entity Generator_sv_unit is
end Generator_sv_unit;
