//****************************************************************************************************  
//*---------------Copyright (c) 2016 C-L-G.FPGA1988.lichangbeiju. All rights reserved-----------------
//
//                   --              It to be define                --
//                   --                    ...                      --
//                   --                    ...                      --
//                   --                    ...                      --
//**************************************************************************************************** 
//File Information
//**************************************************************************************************** 
//File Name      : Monitor.sv 
//Project Name   : azpr_soc_tb
//Description    : the testbench monitor : do some monite and record.
//Github Address : github.com/C-L-G/azpr_soc/trunk/ic/fpga/simulate/tb/Monitor.sv
//License        : Apache-2.0
//**************************************************************************************************** 
//Version Information
//**************************************************************************************************** 
//Create Date    : 2016-12-01 09:00
//First Author   : lichangbeiju
//Last Modify    : 2016-12-01 14:20
//Last Author    : lichangbeiju
//Version Number : 12 commits 
//**************************************************************************************************** 
//Change History(latest change first)
//yyyy.mm.dd - Author - Your log of change
//**************************************************************************************************** 
//2016.12.01 - lichangbeiju - The first version.
//*---------------------------------------------------------------------------------------------------
//File Include : system header file
`include "nettype.h"
`include "global_config.h"
`include "stddef.h"

//File Include : testbench include


`ifndef INC_MONITOR_SV
`define INC_MONITOR_SV
//************************************************************************************************
// 1.Class
//************************************************************************************************

class Monitor;
    //------------------------------------------------------------------------------------------------
    //1.1 Interface define
    //------------------------------------------------------------------------------------------------
    virtual soc_if.iic  iic_if  ;
    
    //------------------------------------------------------------------------------------------------
    //1.2 Class define
    //------------------------------------------------------------------------------------------------   
    

    //------------------------------------------------------------------------------------------------
    //1.3 mailbox define
    //------------------------------------------------------------------------------------------------  
    mailbox             g2d     ;
    mailbox             g2m     ;
    mailbox             d2m     ;
    mailbox             m2s     ;
    

    //------------------------------------------------------------------------------------------------
    //1.4 function and task define
    //------------------------------------------------------------------------------------------------  
    extern function new(virtual soc_if soc_if_i,mailbox d2m_i,m2s_i);
//    extern task recv_data();
    

endclass : Monitor

//************************************************************************************************
//2.Task and function
//************************************************************************************************

//------------------------------------------------------------------------------------------------
//2.1 new function
//------------------------------------------------------------------------------------------------
function Monitor::new(virtual soc_if soc_if_i,mailbox d2m_i,m2s_i);
    this.iic_if = soc_if_i.iic;
    this.d2m    = d2m_i;
    this.m2s    = m2s_i;
endfunction


//------------------------------------------------------------------------------------------------
// 2.2 the send data generator
//------------------------------------------------------------------------------------------------    
//task Monitor::recv_data();

//endtask


`endif
//****************************************************************************************************
//End of Class
//****************************************************************************************************
