library verilog;
use verilog.vl_types.all;
entity Monitor_sv_unit is
end Monitor_sv_unit;
