//****************************************************************************************************  
//*---------------Copyright (c) 2016 C-L-G.FPGA1988.lichangbeiju. All rights reserved-----------------
//
//                   --              It to be define                --
//                   --                    ...                      --
//                   --                    ...                      --
//                   --                    ...                      --
//**************************************************************************************************** 
//File Information
//**************************************************************************************************** 
//File Name      : Scoreboard.sv 
//Project Name   : azpr_soc_tb
//Description    : the testbench scoreboard : compare the result between dut and ref.
//Github Address : github.com/C-L-G/azpr_soc/trunk/ic/fpga/simulate/tb/Scoreboard.sv
//License        : Apache-2.0
//**************************************************************************************************** 
//Version Information
//**************************************************************************************************** 
//Create Date    : 2016-12-01 09:00
//First Author   : lichangbeiju
//Last Modify    : 2016-12-01 14:20
//Last Author    : lichangbeiju
//Version Number : 12 commits 
//**************************************************************************************************** 
//Change History(latest change first)
//yyyy.mm.dd - Author - Your log of change
//**************************************************************************************************** 
//2016.12.02 - lichangbeiju - The first version.
//*---------------------------------------------------------------------------------------------------
//File Include : system header file
`include "nettype.h"
`include "global_config.h"
`include "stddef.h"

//File Include : testbench include


`ifndef INC_SCOREBOARD_SV
`define INC_SCOREBOARD_SV
//************************************************************************************************
// 1.Class
//************************************************************************************************

class Scoreboard;
    //------------------------------------------------------------------------------------------------
    //1.1 Interface define
    //------------------------------------------------------------------------------------------------
    
    //------------------------------------------------------------------------------------------------
    //1.2 Class define
    //------------------------------------------------------------------------------------------------   
    

    //------------------------------------------------------------------------------------------------
    //1.3 mailbox define
    //------------------------------------------------------------------------------------------------  
    mailbox             m2s     ;
    mailbox             g2s     ;
    mailbox             r2s     ;

    

    //------------------------------------------------------------------------------------------------
    //1.4 function and task define
    //------------------------------------------------------------------------------------------------  
    extern function new(mailbox m2s_i,g2s_i);
    extern task comp_run();
    extern task write_read_comp(input bit [07:00] wdata,input bit [07:00] rdata);

endclass : Scoreboard

//************************************************************************************************
//2.Task and function
//************************************************************************************************

//------------------------------------------------------------------------------------------------
//2.1 new function
//------------------------------------------------------------------------------------------------
function Scoreboard::new(mailbox m2s_i,g2s_i);
    this.m2s = m2s_i;
    this.g2s = g2s_i;
endfunction


//------------------------------------------------------------------------------------------------
// 2.2 the send data generator
//------------------------------------------------------------------------------------------------    
task Scoreboard::comp_run();
    logic   [07:00]     m2s_recv    ;
    logic   [07:00]     g2s_recv    ;
    logic               comp_fail   ;
    int                 m2s_num     ;
    int                 g2s_num     ;

    m2s_num     = m2s.num();
    g2s_num     = g2s.num();
    comp_fail   = 0;
    $display("");
    $display("");
    if(m2s_num == g2s_num)
        begin
            for(int i=0;i<g2s_num;i++) begin
                m2s.get(m2s_recv);
                g2s.get(g2s_recv);
                if(g2s_recv == m2s_recv)
                    begin
                        $display("mailbox %0dth data is same : m2s %h = g2s %h.",i,m2s_recv,g2s_recv);
                    end
                else
                    begin
                        comp_fail = 1;
                        $display("mailbox %0dth data is different : the expect data = %h,the read data = %h.",i,g2s_recv,m2s_recv);
                    end
            end
            if(~comp_fail)
                begin
                    $display("//**************************************************************************//");
                    $display("                            Compare success                                   ");
                    $display("//**************************************************************************//");
                end
            else
                begin
                    $display("//**************************************************************************//");
                    $display("                            Compare Fail                                      ");
                    $display("//**************************************************************************//");
                end
        end
    else
        begin
            $display("//**************************************************************************//");
            $display("                            Compare Fail                                      ");
            $display("****The number is different!!!****");
            $display("//**************************************************************************//");

        end
endtask

//------------------------------------------------------------------------------------------------
// 2.3 the write and read data compare
//------------------------------------------------------------------------------------------------    
task Scoreboard::write_read_comp(input bit [07:00] wdata,input bit [07:00] rdata);
    logic           error   ;
    if(wdata != rdata)
        error = 1;
endtask


`endif
//****************************************************************************************************
//End of Class
//****************************************************************************************************
