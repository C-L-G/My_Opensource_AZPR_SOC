//****************************************************************************************************  
//*---------------Copyright (c) 2016 C-L-G.FPGA1988.lichangbeiju. All rights reserved-----------------
//
//                   --              It to be define                --
//                   --                    ...                      --
//                   --                    ...                      --
//                   --                    ...                      --
//**************************************************************************************************** 
//File Information
//**************************************************************************************************** 
//File Name      : Environment.sv 
//Project Name   : azpr_soc_tb
//Description    : the testbench environment.
//Github Address : github.com/C-L-G/azpr_soc/trunk/ic/fpga/simulate/tb/Environment.sv
//License        : Apache-2.0
//**************************************************************************************************** 
//Version Information
//**************************************************************************************************** 
//Create Date    : 2016-12-01 09:00
//First Author   : lichangbeiju
//Last Modify    : 2016-12-01 14:20
//Last Author    : lichangbeiju
//Version Number : 12 commits 
//**************************************************************************************************** 
//Change History(latest change first)
//yyyy.mm.dd - Author - Your log of change
//**************************************************************************************************** 
//2016.12.01 - lichangbeiju - The first version.
//*---------------------------------------------------------------------------------------------------
//File Include : system header file
`include "nettype.h"
`include "global_config.h"
`include "stddef.h"

//File Include : testbench include
`include "Driver.sv"
`include "Generator.sv"
`include "Scoreboard.sv"
`include "Monitor.sv"
//`include "Receiver.sv"
//`include "Reference.sv"

`ifndef INC_ENVIRONMENT_SV
`define INC_ENVIRONMENT_SV
//************************************************************************************************
// 1.Class
//************************************************************************************************

class Environment;
    //------------------------------------------------------------------------------------------------
    //1.1 Interface define
    //------------------------------------------------------------------------------------------------
//    virtual soc_if soc_if       ;
//    virtual soc_if.uart uart_if ;
    
    //------------------------------------------------------------------------------------------------
    //1.2 Class define
    //------------------------------------------------------------------------------------------------   
    Driver              drv     ;
    Generator           gen     ;
    Monitor             mon     ;
    Scoreboard          sb      ;
    

    //------------------------------------------------------------------------------------------------
    //1.3 mailbox define
    //------------------------------------------------------------------------------------------------  
    mailbox             g2d     ;
    mailbox             g2s     ;
    mailbox             m2s     ;
    mailbox             d2m     ;
    

    //------------------------------------------------------------------------------------------------
    //1.4 function and task define
    //------------------------------------------------------------------------------------------------  
    extern function new(virtual soc_if soc_if_i);
    

endclass

//************************************************************************************************
//2.Task and function
//************************************************************************************************

//------------------------------------------------------------------------------------------------
//2.1 new
//------------------------------------------------------------------------------------------------
function Environment::new(virtual soc_if soc_if_i);
//    iic_if.sdo  = 1;
    g2d         = new();
    g2s         = new();
    d2m         = new();
    m2s         = new();
    drv         = new(soc_if_i,g2d,d2m);
    gen         = new(g2d,g2s);
    mon         = new(soc_if_i,d2m,d2m);
    sb          = new(d2m,g2s);
endfunction


//------------------------------------------------------------------------------------------------
// 2.1 the clk generate module
//------------------------------------------------------------------------------------------------    

//------------------------------------------------------------------------------------------------
// 2.2 the interface
//------------------------------------------------------------------------------------------------    

//------------------------------------------------------------------------------------------------
// 2.3 the testcase with interface
//------------------------------------------------------------------------------------------------    

//------------------------------------------------------------------------------------------------
// 2.4 the interface
//------------------------------------------------------------------------------------------------    

//------------------------------------------------------------------------------------------------
// 2.5 the interface
//------------------------------------------------------------------------------------------------    



`endif
//****************************************************************************************************
//End of Class
//****************************************************************************************************
