library verilog;
use verilog.vl_types.all;
entity Environment_sv_unit is
end Environment_sv_unit;
