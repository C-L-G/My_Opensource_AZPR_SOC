library verilog;
use verilog.vl_types.all;
entity Driver_sv_unit is
end Driver_sv_unit;
