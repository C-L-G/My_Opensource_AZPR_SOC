//****************************************************************************************************  
//*---------------Copyright (c) 2016 C-L-G.FPGA1988.lichangbeiju. All rights reserved-----------------
//
//                   --              It to be define                --
//                   --                    ...                      --
//                   --                    ...                      --
//                   --                    ...                      --
//**************************************************************************************************** 
//File Information
//**************************************************************************************************** 
//File Name      : Generator.sv 
//Project Name   : azpr_soc_tb
//Description    : the testbench generator : gen the data and send it to the drv or scoreboard.
//Github Address : github.com/C-L-G/azpr_soc/trunk/ic/fpga/simulate/tb/Generator.sv
//License        : Apache-2.0
//**************************************************************************************************** 
//Version Information
//**************************************************************************************************** 
//Create Date    : 2016-12-01 09:00
//First Author   : lichangbeiju
//Last Modify    : 2016-12-01 14:20
//Last Author    : lichangbeiju
//Version Number : 12 commits 
//**************************************************************************************************** 
//Change History(latest change first)
//yyyy.mm.dd - Author - Your log of change
//**************************************************************************************************** 
//2016.12.01 - lichangbeiju - The first version.
//*---------------------------------------------------------------------------------------------------
//File Include : system header file
`include "nettype.h"
`include "global_config.h"
`include "stddef.h"

//File Include : testbench include


`ifndef INC_GENERATOR_SV
`define INC_GENERATOR_SV
//************************************************************************************************
// 1.Class
//************************************************************************************************

class Generator;
    //------------------------------------------------------------------------------------------------
    //1.1 Interface define
    //------------------------------------------------------------------------------------------------
    
    //------------------------------------------------------------------------------------------------
    //1.2 Class define
    //------------------------------------------------------------------------------------------------   
    

    //------------------------------------------------------------------------------------------------
    //1.3 mailbox define
    //------------------------------------------------------------------------------------------------  
    mailbox             g2d     ;
    mailbox             g2s     ;
    

    //------------------------------------------------------------------------------------------------
    //1.4 function and task define
    //------------------------------------------------------------------------------------------------  
    extern function new(mailbox g2d_i,g2s_i);
    extern task send_data_gen(input bit [07:00] data_start,input bit [15:00] len);
    extern task chk_data_gen(input bit data_same_en,input bit [07:00] data_start,input bit [15:00] len);
    

endclass : Generator

//************************************************************************************************
//2.Task and function
//************************************************************************************************

//------------------------------------------------------------------------------------------------
//2.1 new function
//------------------------------------------------------------------------------------------------
function Generator::new(mailbox g2d_i,g2s_i);
    this.g2d = g2d_i;
    this.g2s = g2s_i;
endfunction


//------------------------------------------------------------------------------------------------
// 2.2 the send data generator
//------------------------------------------------------------------------------------------------    
task Generator::send_data_gen(input bit [07:00] data_start,input bit [15:00] len);
    logic   [07:00]     data = 0    ;
    data     = data_start;
    for(int i = 0;i < len;i++) begin
        g2d.put(data)       ;
        data = data + 1'b1  ;
    end
endtask

//------------------------------------------------------------------------------------------------
// 2.3 the check data generator
//------------------------------------------------------------------------------------------------    
task Generator::chk_data_gen(input bit data_same_en,input bit [07:00] data_start,input bit [15:00] len);
    logic   [07:00]     data = 0    ;
    data    = data_start;
    for(int i = 0;i < len;i++) begin
        g2s.put(data);
        if(~data_same_en)
            data = data + 1'b1;
        else
            data = data;
    end
endtask


`endif
//****************************************************************************************************
//End of Class
//****************************************************************************************************
