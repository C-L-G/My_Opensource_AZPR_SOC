//****************************************************************************************************  
//*---------------Copyright (c) 2016 C-L-G.FPGA1988.lichangbeiju. All rights reserved-----------------
//
//                   --              It to be define                --
//                   --                    ...                      --
//                   --                    ...                      --
//                   --                    ...                      --
//**************************************************************************************************** 
//File Information
//**************************************************************************************************** 
//File Name      : Testbench.sv 
//Project Name   : azpr_soc
//Description    : the fpga testbench top of the chip.
//Github Address : github.com/C-L-G/azpr_soc/trunk/ic/fpga/simulate/tb/Testbench.sv
//License        : Apache-2.0
//**************************************************************************************************** 
//Version Information
//**************************************************************************************************** 
//Create Date    : 2016-12-01 09:00
//First Author   : lichangbeiju
//Last Modify    : 2016-12-01 14:20
//Last Author    : lichangbeiju
//Version Number : 12 commits 
//**************************************************************************************************** 
//Change History(latest change first)
//yyyy.mm.dd - Author - Your log of change
//**************************************************************************************************** 
//2016.12.01 - lichangbeiju - The first version.
//*---------------------------------------------------------------------------------------------------
//File Include : system header file
`include "nettype.h"
`include "global_config.h"
`include "stddef.h"

module clock_reset(
    output  bit         system_clock    ,
    output  bit         reset


);
    //************************************************************************************************
    // 1.Parameter and constant define
    //***********************************************************************************************
    localparam CLOCK_LOW_TIME   = 10    ;
    localparam CLOCK_HIGH_TIME  = 10    ;
    
    //************************************************************************************************
    // 2.Register and wire declaration
    //************************************************************************************************
    //------------------------------------------------------------------------------------------------
    // 2.1 the output reg
    //------------------------------------------------------------------------------------------------   
    logic                   sda_m2s     ;
    logic   [00:00]         sda_s2m     ;
    logic                   scl         ;
    logic                   clk         ;
    //------------------------------------------------------------------------------------------------
    // 2.2 the internal reg
    //------------------------------------------------------------------------------------------------  
    
    logic                   sample_flag ;//bus inteface state
    int                     fp_eeprom   ;//
    bit                     vect_clk    ;//vector clock


    reg                     ck_en       ;
    //------------------------------------------------------------------------------------------------
    // 2.x the test logic
    //------------------------------------------------------------------------------------------------

    //************************************************************************************************
    // 3.Main code
    //************************************************************************************************

    //------------------------------------------------------------------------------------------------
    // 3.1 the sdf annotate 
    //------------------------------------------------------------------------------------------------
    initial begin
        system_clock = 1'b0 ;
        ck_en        = 1'b1 ;
    end

    initial begin
        reset = `RESET_ENABLE   ;
        #100;
        reset = `RESET_DISABLE  ;

    end


    //------------------------------------------------------------------------------------------------
    // 3.2 the signal assignment
    //------------------------------------------------------------------------------------------------
    task run(int reset_hold = 4,int l_period = CLOCK_LOW_TIME,int h_period = CLOCK_HIGH_TIME,int count=0);
        system_clock = 0;
        for(int clk_i=0;(clk_i < count  || count == 0);clk_i++)
            if(ck_en)
                #l_period;
                    system_clock = ~system_clock;
                #h_period;
                    system_clock = ~system_clock;
            else
                system_clock = 1'b0;
    endtask
    //------------------------------------------------------------------------------------------------
    // 3.4 the hsim vector generate
    //------------------------------------------------------------------------------------------------
    `ifdef hsim
        initial begin : VECTOR_GEN_INIT
            fp_eeprom = $fopen("./hsim.vec","w+");
            
            $fdisplay(fp_eeprom,"radix  1       1       1       1   \n");
            $fdisplay(fp_eeprom,"io     i       i       i       i   \n");
            $fdisplay(fp_eeprom,"vname  pad1    pad3    pad5    pad6\n");

            $fdisplay(fp_eeprom,"period 10 ");
            $fdisplay(fp_eeprom,"TUNIT  1ns");
            $fdisplay(fp_eeprom,"vih    simvih");
            $fdisplay(fp_eeprom,"tskip");
            $fdisplay(fp_eeprom,"\n");
        end
        
        initial begin
            vect_clk    = 1'b0;
        end
        always begin
            #10 vect_clk = ~vect_clk;
        end 
        
        always @(posedge vect_clk) begin : VECTOR_GEN_SAMPLE
            if(sample_flag)
                $fdisplay(fp_eeprom,"%10d   %h  %h  %h  %h",
                $time,test_top.pad1,test_top.pad3,test_top.pad5,test_top.pad6);
        end
    `endif

    //************************************************************************************************
    // 4.Sub module instantiation
    //************************************************************************************************
    //------------------------------------------------------------------------------------------------
    // 4.1 the clk generate module
    //------------------------------------------------------------------------------------------------    
    azpr_clock_reset cr(.*);

    //------------------------------------------------------------------------------------------------
    // 4.2 the interface
    //------------------------------------------------------------------------------------------------    
    soc_if soc_if(system_clock);
    
    //------------------------------------------------------------------------------------------------
    // 4.3 the testcase with interface
    //------------------------------------------------------------------------------------------------    
    testcase tc(soc_if);
    
    //------------------------------------------------------------------------------------------------
    // 4.4 the interface
    //------------------------------------------------------------------------------------------------    
    gt5232_chip_top dut(.*);

    //------------------------------------------------------------------------------------------------
    // 4.5 the interface
    //------------------------------------------------------------------------------------------------    




endmodule    
//****************************************************************************************************
//End of Mopdule
//****************************************************************************************************
