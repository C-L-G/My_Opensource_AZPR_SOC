library verilog;
use verilog.vl_types.all;
entity Scoreboard_sv_unit is
end Scoreboard_sv_unit;
