library verilog;
use verilog.vl_types.all;
entity Testbench is
end Testbench;
