//****************************************************************************************************  
//*---------------Copyright (c) 2016 C-L-G.FPGA1988.lichangbeiju. All rights reserved-----------------
//
//                   --              It to be define                --
//                   --                    ...                      --
//                   --                    ...                      --
//                   --                    ...                      --
//**************************************************************************************************** 
//File Information
//**************************************************************************************************** 
//File Name      : clock_reset.sv 
//Project Name   : azpr_soc
//Description    : the fpga testbench clock reset.
//Github Address : github.com/C-L-G/azpr_soc/trunk/ic/fpga/simulate/tb/Testbench.sv
//License        : Apache-2.0
//**************************************************************************************************** 
//Version Information
//**************************************************************************************************** 
//Create Date    : 2016-12-01 09:00
//First Author   : lichangbeiju
//Last Modify    : 2016-12-23 14:20
//Last Author    : lichangbeiju
//Version Number : 12 commits 
//**************************************************************************************************** 
//Change History(latest change first)
//yyyy.mm.dd - Author - Your log of change
//**************************************************************************************************** 
//2016.12.23 - lichangbeiju - Add the cr.run task.
//2016.12.01 - lichangbeiju - The first version.
//*---------------------------------------------------------------------------------------------------
//File Include : system header file
`include "nettype.h"
`include "global_config.h"
`include "stddef.h"

module clock_reset(
    output  bit         system_clock    ,
    output  bit         reset


);
    //************************************************************************************************
    // 1.Parameter and constant define
    //***********************************************************************************************
    localparam CLOCK_LOW_TIME   = 10    ;
    localparam CLOCK_HIGH_TIME  = 10    ;
    
    //************************************************************************************************
    // 2.Register and wire declaration
    //************************************************************************************************
    //------------------------------------------------------------------------------------------------
    // 2.1 the output reg
    //------------------------------------------------------------------------------------------------   
    reg                     ck_en       ;

    //------------------------------------------------------------------------------------------------
    // 2.x the test logic
    //------------------------------------------------------------------------------------------------

    //************************************************************************************************
    // 3.Main code
    //************************************************************************************************

    //------------------------------------------------------------------------------------------------
    // 3.1 the sdf annotate 
    //------------------------------------------------------------------------------------------------
    initial begin
        system_clock = 1'b0 ;
        ck_en        = 1'b1 ;
    end

    initial begin
        reset = `RESET_ENABLE   ;
        #100;
        reset = `RESET_DISABLE  ;

    end

    //------------------------------------------------------------------------------------------------
    // 3.2 the signal assignment
    //------------------------------------------------------------------------------------------------
    task run(int reset_hold = 4,int l_period = CLOCK_LOW_TIME,int h_period = CLOCK_HIGH_TIME,int count=0);
        system_clock = 0;
        for(int clk_i=0;(clk_i < count  || count == 0);clk_i++)
            if(ck_en) begin
                #l_period;
                    system_clock = ~system_clock;
                #h_period;
                    system_clock = ~system_clock;
			end
            else
                system_clock = 1'b0;
    endtask
    //------------------------------------------------------------------------------------------------
    // 3.4 the hsim vector generate
    //------------------------------------------------------------------------------------------------

    //************************************************************************************************
    // 4.Sub module instantiation
    //************************************************************************************************
    //------------------------------------------------------------------------------------------------
    // 4.1 the clk generate module
    //------------------------------------------------------------------------------------------------    

endmodule    
//****************************************************************************************************
//End of Mopdule
//****************************************************************************************************
